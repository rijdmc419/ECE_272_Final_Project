module decoder #(parameter N = 8, M = 10)(input logic [N-1:0] in,
														 output logic [16:0] y);
		
			//need a 17 bit output b/c max number for A half flat under A 440 needs 17 bits
			always_comb	
			case(in)
		 
			28: y = 113636.3636; //A
			27: y = 107259.3101; //S
			35: y = 101239.1674; //D
			/*43: y = 95556.6173; //F
			52: y = 90192.47073; //G
			51: y = 85131.01663; //H
			59: y = 80353.55564; //J
			66: y = 75843.76185; //K
			75: y = 71586.06076; //L
			76: y = 67568.48066; //;
			82: y = 63776.32368; //'
			90: y = 60196.72289; //enter
			
			21: y = 116967.2726; //Q
			29: y = 110402.0844; //W
			36: y = 104205.7438; //E
			45: y = 98356.46349; //R
			44: y = 92836.71878; //T
			53: y = 87627.05924; //Y
			60: y = 82712.98594; //U
			67: y = 78066.45016; //I
			68: y = 73684.36565; //O
			77: y = 69548.7676; //P
			84: y = 65645.22694; //[
			91: y = 61960.93982; //]
			
			18: y = 110402.0844; //Left shift
			26: y = 104205.7438; //Z
			34: y = 98356.46349; //X
			33: y = 92836.71878; //C
			42: y = 87627.05924; //V
			50: y = 82712.98594; //B
			49: y = 78066.45016; //N
			58: y = 73684.36565; //M
			65: y = 69548.7676; //,
			73: y = 65645.22694; //.
			74: y = 61960.93982; // /
			89: y = 58483.63628; //right shift
			*/
			default: y=0;
			
			endcase
			
			
			
endmodule